package cfg;
	bit clk_100khz; 
endpackage
