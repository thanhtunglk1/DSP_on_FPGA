module TWI_FSM_master #(
    parameter SIZE_CMD = 3
)(
    input logic                     i_clk   ,
    input logic                     i_rst_n ,
    input logic                     i_TWIEN ,
    input logic [SIZE_CMD-1:0]      i_cmd   ,
     
);

endmodule

