`include "design.sv"
`include "dut_interface.sv"
`include "trans1.svh"
`include "tr_sequence.svh"
`include "tb_sequencer.svh"
`include "tb_driver.svh"
`include "tb_monitor.svh"
`include "tb_scoreboard.svh"
`include "tb_agent.svh"
`include "tb_environment.svh"
`include "base_test.svh"
`include "sanity_test.svh"
`include "full_memory_test.svh"
